`timescale 1ns / 1ps

//top module test bench




module tb_top_module();

    parameter DSIZE = 8; // Data bus size
    parameter ASIZE = 4; // Address bus size
    parameter DEPTH = 1 << ASIZE; // Depth of the FIFO memory

    reg [DSIZE-1:0] wdata;   // Input data
    wire [DSIZE-1:0] rdata;  // Output data
    wire wfull, rempty, walmost_full, ralmost_empty;      // Write full and read empty signals
    reg winc, rinc, wclk, rclk, wrst_n, rrst_n; // Write and read signals
//    wire [3:0] waddr, raddr;

    top_module #(.n(ASIZE), .DATA(DSIZE), .DEPTH(ASIZE)) FIFO (
        .wclk(wclk),
        .rclk(rclk),
        .wrst_n(wrst_n),
        .rrst_n(rrst_n),
        .winc(winc),
        .rinc(rinc),
        .wdata(wdata),

        .rdata(rdata),
        .wfull(wfull),
        .rempty(rempty),
        .walmost_full(walmost_full),
        .ralmost_empty(ralmost_empty)
//        .w_bptr(waddr), .r_bptr(raddr)
    );

    integer i=0;
    integer seed = 1;

    // Read and write clock in loop
    always #5 wclk = ~wclk;    // faster writing
    always #10 rclk = ~rclk;   // slower reading
    
    initial begin
        // Initialize all signals
        wclk = 0;
        rclk = 0;
        wrst_n = 0;     // Active low reset
        rrst_n = 0;     // Active low reset
        winc = 0;
        rinc = 0;
        wdata = 0;

        // Reset the FIFO
        #100 wrst_n = 0; rrst_n = 0;
        #40 wrst_n = 1; rrst_n = 1;

        // TEST CASE 1: Write data and read it back
//         rinc = 1;
//         for (i = 0; i < 40; i = i + 1) begin
//             wdata = $random(seed) % 256;
//             winc = 1;
//             #10;
//             winc = 0;
//             #10;
//         end

        // TEST CASE 2: Write data to make FIFO full and try to write more data
//        rinc = 0;
//        winc = 1;
//        for (i = 0; i < DEPTH + 3; i = i + 1) begin
//            wdata = $random(seed) % 256;
//            #10;
//        end

//        #30

        // TEST CASE 3: Read data from empty FIFO and try to read more data
//        winc = 0;
//        rinc = 1;
//        for (i = 0; i < DEPTH + 3; i = i + 1) begin
//            #20;
//        end

        // TEST CASE 4: Write 2 data and read 1 data
         // for (i = 0; i < 20; i = i + 1) begin
         //     wdata = $random(seed) % 256;
         //     winc = 1;
         //     #10;
         //     wdata = $random(seed) % 256;
         //     #10;
         //     winc=0; rinc=1;
         //     #20
         //     rinc=0;
         // end

        // TEST CASE 5: Write until fifo become full and then read until fifo become empty
        rinc = 0;
        winc = 1;
        for (i = 0; i < DEPTH + 4; i = i + 1) begin
            wdata = $random(seed) % 256;
            #10;
        end
        winc = 0;
        #30
        rinc = 1;
        for (i = 0; i < DEPTH + 3; i = i + 1) begin
            #20;
        end

        $stop;
    end

endmodule
